module and_gate(input a, b, output x);

and and1 (x, a, b);

endmodule
