module FirstPain (input a, b, output s);

and and1 (s, a, b);

end module;

